import "DPI-C" function int serial_tick
(
    input  bit     serial_out_valid,
    output bit     serial_out_ready,
    input  int     serial_out_bits,

    output bit     serial_in_valid,
    input  bit     serial_in_ready,
    output int     serial_in_bits,

    input int      nchannels,
    input longint  mem_size,
    input int      word_bytes,
    input int      line_bytes,
    input int      id_bits
);

module SimSerial #(
    parameter SERIAL_WIDTH = 32,
              NUM_CHANNELS = 1,
              MEM_SIZE = 1000 * 1000 * 1000,
              WORD_BYTES = 8,
              LINE_BYTES = 64,
              ID_BITS = 5)
(
    input                     clock,
    input                     reset,
    input                     serial_out_valid,
    output                    serial_out_ready,
    input  [SERIAL_WIDTH-1:0] serial_out_bits,

    output                    serial_in_valid,
    input                     serial_in_ready,
    output [SERIAL_WIDTH-1:0] serial_in_bits,

    output                     exit
);

    bit __in_valid;
    bit __out_ready;
    int __in_bits;
    int __exit;

    reg __in_valid_reg;
    reg __out_ready_reg;
    reg [31:0] __in_bits_reg;
    reg __exit_reg;

    assign serial_in_valid  = __in_valid_reg;
    assign serial_in_bits   = __in_bits_reg;
    assign serial_out_ready = __out_ready_reg;
    assign exit = __exit_reg;

    // Evaluate the signals on the positive edge
    always @(posedge clock) begin
        if (reset) begin
            __in_valid = 0;
            __out_ready = 0;
            __exit = 0;

            __in_valid_reg <= 0;
            __in_bits_reg <= 0;
            __out_ready_reg <= 0;
            __exit_reg <= 0;
        end else begin
            __exit = serial_tick(
                serial_out_valid,
                __out_ready,
                serial_out_bits,
                __in_valid,
                serial_in_ready,
                __in_bits,
                NUM_CHANNELS,
                MEM_SIZE,
                WORD_BYTES,
                LINE_BYTES,
                ID_BITS
            );

            __out_ready_reg <= __out_ready;
            __in_valid_reg  <= __in_valid;
            __in_bits_reg   <= __in_bits;
            __exit_reg <= __exit[0];
        end
    end

endmodule
